module freeList # (

) (

);