module RAT # (
    parameter CORE_WIDTH = 2
) (

);


endmodule
