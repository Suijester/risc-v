// decode-rename pipeline buffer