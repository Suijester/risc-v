module controlUnit (
    input logic 
);

endmodule